"1+1";