for(let i=1;i<5;i++) g=2 ;
do   document.write(" bye 2 "); while(i!=5)