{a:5, "k":"yanny", c:2+3*8 || 3+3, [9+9*2]:"esteban", y:[2,3,4], f:[]};