"a" | upper