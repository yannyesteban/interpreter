yanny { @home } esteban {{ @a }} siempre {{ @b }}

yanny {@name} r: {@age} nothing {@k.b.1 | upper}
{@price | digits:2 | format} {@birth | date}
{@_DATE_} {@_TIME_}