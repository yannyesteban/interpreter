let name = {a:2}; name.a | upper