yanny {@name} r: {@age} nothing {@k.b.1 | upper}