yanny {@name} r: {@age} nothing