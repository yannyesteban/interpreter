func a(){return 1};
a()