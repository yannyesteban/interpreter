{a:5};