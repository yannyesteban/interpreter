{: 2+2 :}