a + c ** d ** YAnny;