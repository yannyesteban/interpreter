if(1+2){2+2}