a:={b:1};
a.b++;
a.b