a("p");