func x(a){
    a+36
}

x(9)