a:=5;
a;
a++
a