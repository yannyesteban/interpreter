"yanny";
let name = {
    "a": {
        "name": "yanny",
        "last": "jimenez"
    }
};
name.a.last | upper;