math.cos(45)