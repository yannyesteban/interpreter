g=2;if(a>2)l=9;