let name = "yanny"; name | upper