"yanny";
let name = {a:{name:"yanny",last:"nuñez"}};
name.a.last | upper;