{if(a>1)d=9}