++5;